--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   17:40:58 05/14/2019
-- Design Name:   
-- Module Name:   /home/calvillo/Bureau/Compilateur/VHDL/Processeur/MemoireTB.vhd
-- Project Name:  Processeur
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: MemoireDonnees
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY MemoireTB IS
END MemoireTB;
 
ARCHITECTURE behavior OF MemoireTB IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT MemoireDonnees
    PORT(
         addr : IN  std_logic_vector(3 downto 0);
         Input : IN  std_logic_vector(15 downto 0);
         RW : IN  std_logic;
         RST : IN  std_logic;
         CLK : IN  std_logic;
         Output : OUT  std_logic_vector(15 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal addr : std_logic_vector(3 downto 0) := (others => '0');
   signal Input : std_logic_vector(15 downto 0) := (others => '0');
   signal RW : std_logic := '0';
   signal RST : std_logic := '0';
   signal CLK : std_logic := '0';

 	--Outputs
   signal Output : std_logic_vector(15 downto 0);

   -- Clock period definitions
   constant CLK_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: MemoireDonnees PORT MAP (
          addr => addr,
          Input => Input,
          RW => RW,
          RST => RST,
          CLK => CLK,
          Output => Output
        );

   -- Clock process definitions
   CLK_process :process
   begin
		CLK <= '0';
		wait for CLK_period/2;
		CLK <= '1';
		wait for CLK_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      RST <= '1';
		wait for 100 ns;	
		RST <= '0';
		
      wait for CLK_period*10;
		addr <= x"0";
		input <= x"FFFF";
		RW <= '0';
		wait for CLK_period*10;
      
		addr <= x"0";
		input <= x"0001";
		RW <= '1';
		wait for CLK_period*10;
      RST <= '1';
		wait for CLK_period*10;
      
		
		-- insert stimulus here 

      wait;
   end process;

END;
